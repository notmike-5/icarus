// helpful encoders

module priority_encode #(parameter N = 255)
  (
    input		       en,
    input [N-1:0]	       n,
    output reg [$clog2(N)-1:0] i
   );

  always @(en, n)
    assign i = (!en) ? 8'bzzzzzzzz :
	       (n[254]) ? 8'd254 : 
	       (n[253]) ? 8'd253 :
	       (n[252]) ? 8'd252 : 
	       (n[251]) ? 8'd251 :
	       (n[250]) ? 8'd250 :
	       (n[249]) ? 8'd249 :
	       (n[248]) ? 8'd248 :
	       (n[247]) ? 8'd247 :
	       (n[246]) ? 8'd246 :
	       (n[245]) ? 8'd245 :
	       (n[244]) ? 8'd244 :
	       (n[243]) ? 8'd243 :
	       (n[242]) ? 8'd242 :
	       (n[241]) ? 8'd241 :
	       (n[240]) ? 8'd240 :
	       (n[239]) ? 8'd239 :
	       (n[238]) ? 8'd238 :
	       (n[237]) ? 8'd237 :
	       (n[236]) ? 8'd236 :
	       (n[235]) ? 8'd235 :
	       (n[234]) ? 8'd234 :
	       (n[233]) ? 8'd233 :
	       (n[232]) ? 8'd232 :
	       (n[231]) ? 8'd231 :
	       (n[230]) ? 8'd230 :
	       (n[229]) ? 8'd229 :
	       (n[228]) ? 8'd228 :
	       (n[227]) ? 8'd227 :
	       (n[226]) ? 8'd226 :
	       (n[225]) ? 8'd225 :
	       (n[224]) ? 8'd224 :
	       (n[223]) ? 8'd223 :
	       (n[222]) ? 8'd222 :
	       (n[221]) ? 8'd221 :
	       (n[220]) ? 8'd220 :
	       (n[219]) ? 8'd219 :
	       (n[218]) ? 8'd218 :
	       (n[217]) ? 8'd217 :
	       (n[216]) ? 8'd216 :
	       (n[215]) ? 8'd215 :
	       (n[214]) ? 8'd214 :
	       (n[213]) ? 8'd213 :
	       (n[212]) ? 8'd212 :
	       (n[211]) ? 8'd211 :
	       (n[210]) ? 8'd210 :
	       (n[209]) ? 8'd209 :
	       (n[208]) ? 8'd208 :
	       (n[207]) ? 8'd207 :
	       (n[206]) ? 8'd206 :
	       (n[205]) ? 8'd205 :
	       (n[204]) ? 8'd204 :
	       (n[203]) ? 8'd203 :
	       (n[202]) ? 8'd202 :
	       (n[201]) ? 8'd201 :
	       (n[200]) ? 8'd200 :
	       (n[199]) ? 8'd199 :
	       (n[198]) ? 8'd198 :
	       (n[197]) ? 8'd197 :
	       (n[196]) ? 8'd196 :
	       (n[195]) ? 8'd195 :
	       (n[194]) ? 8'd194 :
	       (n[193]) ? 8'd193 :
	       (n[192]) ? 8'd192 :
	       (n[191]) ? 8'd191 :
	       (n[190]) ? 8'd190 :
	       (n[189]) ? 8'd189 :
	       (n[188]) ? 8'd188 :
	       (n[187]) ? 8'd187 :
	       (n[186]) ? 8'd186 :
	       (n[185]) ? 8'd185 :
	       (n[184]) ? 8'd184 :
	       (n[183]) ? 8'd183 :
	       (n[182]) ? 8'd182 :
	       (n[181]) ? 8'd181 :
	       (n[180]) ? 8'd180 :
	       (n[179]) ? 8'd179 :
	       (n[178]) ? 8'd178 :
	       (n[177]) ? 8'd177 :
	       (n[176]) ? 8'd176 :
	       (n[175]) ? 8'd175 :
	       (n[174]) ? 8'd174 :
	       (n[173]) ? 8'd173 :
	       (n[172]) ? 8'd172 :
	       (n[171]) ? 8'd171 :
	       (n[170]) ? 8'd170 :
	       (n[169]) ? 8'd169 :
	       (n[168]) ? 8'd168 :
	       (n[167]) ? 8'd167 :
	       (n[166]) ? 8'd166 :
	       (n[165]) ? 8'd165 :
	       (n[164]) ? 8'd164 :
	       (n[163]) ? 8'd163 :
	       (n[162]) ? 8'd162 :
	       (n[161]) ? 8'd161 :
	       (n[160]) ? 8'd160 :
	       (n[159]) ? 8'd159 :
	       (n[158]) ? 8'd158 :
	       (n[157]) ? 8'd157 :
	       (n[156]) ? 8'd156 :
	       (n[155]) ? 8'd155 :
	       (n[154]) ? 8'd154 :
	       (n[153]) ? 8'd153 :
	       (n[152]) ? 8'd152 :
	       (n[151]) ? 8'd151 :
	       (n[150]) ? 8'd150 :
	       (n[149]) ? 8'd149 :
	       (n[148]) ? 8'd148 :
	       (n[147]) ? 8'd147 :
	       (n[146]) ? 8'd146 :
	       (n[145]) ? 8'd145 :
	       (n[144]) ? 8'd144 :
	       (n[143]) ? 8'd143 :
	       (n[142]) ? 8'd142 :
	       (n[141]) ? 8'd141 :
	       (n[140]) ? 8'd140 :
	       (n[139]) ? 8'd139 :
	       (n[138]) ? 8'd138 :
	       (n[137]) ? 8'd137 :
	       (n[136]) ? 8'd136 :
	       (n[135]) ? 8'd135 :
	       (n[134]) ? 8'd134 :
	       (n[133]) ? 8'd133 :
	       (n[132]) ? 8'd132 :
	       (n[131]) ? 8'd131 :
	       (n[130]) ? 8'd130 :
	       (n[129]) ? 8'd129 :
	       (n[128]) ? 8'd128 :
	       (n[127]) ? 8'd127 :
	       (n[126]) ? 8'd126 :
	       (n[125]) ? 8'd125 :
	       (n[124]) ? 8'd124 :
	       (n[123]) ? 8'd123 :
	       (n[122]) ? 8'd122 :
	       (n[121]) ? 8'd121 :
	       (n[120]) ? 8'd120 :
	       (n[119]) ? 8'd119 :
	       (n[118]) ? 8'd118 :
	       (n[117]) ? 8'd117 :
	       (n[116]) ? 8'd116 :
	       (n[115]) ? 8'd115 :
	       (n[114]) ? 8'd114 :
	       (n[113]) ? 8'd113 :
	       (n[112]) ? 8'd112 :
	       (n[111]) ? 8'd111 :
	       (n[110]) ? 8'd110 :
	       (n[109]) ? 8'd109 :
	       (n[108]) ? 8'd108 :
	       (n[107]) ? 8'd107 :
	       (n[106]) ? 8'd106 :
	       (n[105]) ? 8'd105 :
	       (n[104]) ? 8'd104 :
	       (n[103]) ? 8'd103 :
	       (n[102]) ? 8'd102 :
	       (n[101]) ? 8'd101 :
	       (n[100]) ? 8'd100 :
	       (n[99]) ? 8'd99 :
	       (n[98]) ? 8'd98 :
	       (n[97]) ? 8'd97 :
	       (n[96]) ? 8'd96 :
	       (n[95]) ? 8'd95 :
	       (n[94]) ? 8'd94 :
	       (n[93]) ? 8'd93 :
	       (n[92]) ? 8'd92 :
	       (n[91]) ? 8'd91 :
	       (n[90]) ? 8'd90 :
	       (n[89]) ? 8'd89 :
	       (n[88]) ? 8'd88 :
	       (n[87]) ? 8'd87 :
	       (n[86]) ? 8'd86 :
	       (n[85]) ? 8'd85 :
	       (n[84]) ? 8'd84 :
	       (n[83]) ? 8'd83 :
	       (n[82]) ? 8'd82 :
	       (n[81]) ? 8'd81 :
	       (n[80]) ? 8'd80 :
	       (n[79]) ? 8'd79 :
	       (n[78]) ? 8'd78 :
	       (n[77]) ? 8'd77 :
	       (n[76]) ? 8'd76 :
	       (n[75]) ? 8'd75 :
	       (n[74]) ? 8'd74 :
	       (n[73]) ? 8'd73 :
	       (n[72]) ? 8'd72 :
	       (n[71]) ? 8'd71 :
	       (n[70]) ? 8'd70 :
	       (n[69]) ? 8'd69 :
	       (n[68]) ? 8'd68 :
	       (n[67]) ? 8'd67 :
	       (n[66]) ? 8'd66 :
	       (n[65]) ? 8'd65 :
	       (n[64]) ? 8'd64 :
	       (n[63]) ? 8'd63 :
	       (n[62]) ? 8'd62 :
	       (n[61]) ? 8'd61 :
	       (n[60]) ? 8'd60 :
	       (n[59]) ? 8'd59 :
	       (n[58]) ? 8'd58 :
	       (n[57]) ? 8'd57 :
	       (n[56]) ? 8'd56 :
	       (n[55]) ? 8'd55 :
	       (n[54]) ? 8'd54 :
	       (n[53]) ? 8'd53 :
	       (n[52]) ? 8'd52 :
	       (n[51]) ? 8'd51 :
	       (n[50]) ? 8'd50 :
	       (n[49]) ? 8'd49 :
	       (n[48]) ? 8'd48 :
	       (n[47]) ? 8'd47 :
	       (n[46]) ? 8'd46 :
	       (n[45]) ? 8'd45 :
	       (n[44]) ? 8'd44 :
	       (n[43]) ? 8'd43 :
	       (n[42]) ? 8'd42 :
	       (n[41]) ? 8'd41 :
	       (n[40]) ? 8'd40 :
	       (n[39]) ? 8'd39 :
	       (n[38]) ? 8'd38 :
	       (n[37]) ? 8'd37 :
	       (n[36]) ? 8'd36 :
	       (n[35]) ? 8'd35 :
	       (n[34]) ? 8'd34 :
	       (n[33]) ? 8'd33 :
	       (n[32]) ? 8'd32 :
	       (n[31]) ? 8'd31 :
	       (n[30]) ? 8'd30 :
	       (n[29]) ? 8'd29 :
	       (n[28]) ? 8'd28 :
	       (n[27]) ? 8'd27 :
	       (n[26]) ? 8'd26 :
	       (n[25]) ? 8'd25 :
	       (n[24]) ? 8'd24 :
	       (n[23]) ? 8'd23 :
	       (n[22]) ? 8'd22 :
	       (n[21]) ? 8'd21 :
	       (n[20]) ? 8'd20 :
	       (n[19]) ? 8'd19 :
	       (n[18]) ? 8'd18 :
	       (n[17]) ? 8'd17 :
	       (n[16]) ? 8'd16 :
	       (n[15]) ? 8'd15 :
	       (n[14]) ? 8'd14 :
	       (n[13]) ? 8'd13 :
	       (n[12]) ? 8'd12 :
	       (n[11]) ? 8'd11 :
	       (n[10]) ? 8'd10 :
	       (n[9]) ? 8'd9 :
	       (n[8]) ? 8'd8 :
	       (n[7]) ? 8'd7 :
	       (n[6]) ? 8'd6 :
	       (n[5]) ? 8'd5 :
	       (n[4]) ? 8'd4 :
	       (n[3]) ? 8'd3 :
	       (n[2]) ? 8'd2 :
	       (n[1]) ? 8'd1 : 8'd0;
endmodule
